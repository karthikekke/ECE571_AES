    Mac OS X            	   2  �     �                                    ATTR����  �     �                      com.apple.TextEncoding          com.apple.lastuseddate#PS      '   �  7com.apple.metadata:kMDLabel_noud5bnoeftpfftpczfkpu3kde   utf-8;134217984��ge    ɗ�    �]�S�Z`���9s�\/��E�Xy{]k��}"#C�r��N�L����u2-���$�DYGJ�����P~���RT�
lB}˥�u��q��3RT�)��;�
�4ϫ���+.�w�fw��2��/l��hUг�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               This resource fork intentionally left blank                                                                                                                                                                                                                            ��